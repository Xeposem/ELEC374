library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity encoder32to5 is port(
		input : in std_logic_vector(31 downto 0);
		output: out std_logic_vector(4 downto 0)
);
end entity encoder32to5;

architecture behav of encoder32to5 is
begin
output <= 	  "00000" when (input = "00000000000000000000000000000001")
			else "00001" when (input = "00000000000000000000000000000010")
			else "00010" when (input = "00000000000000000000000000000100")
			else "00011" when (input = "00000000000000000000000000001000")
			else "00100" when (input = "00000000000000000000000000010000")
			else "00101" when (input = "00000000000000000000000000100000")
			else "00110" when (input = "00000000000000000000000001000000")
			else "00111" when (input = "00000000000000000000000010000000")
			else "01000" when (input = "00000000000000000000000100000000")
			else "01001" when (input = "00000000000000000000001000000000")
			else "01010" when (input = "00000000000000000000010000000000")
			else "01011" when (input = "00000000000000000000100000000000")
			else "01100" when (input = "00000000000000000001000000000000")
			else "01101" when (input = "00000000000000000010000000000000")
			else "01110" when (input = "00000000000000000100000000000000")
			else "01111" when (input = "00000000000000001000000000000000")
			else "10000" when (input = "00000000000000010000000000000000")
			else "10001" when (input = "00000000000000100000000000000000")
			else "10010" when (input = "00000000000001000000000000000000")
			else "10011" when (input = "00000000000010000000000000000000")
			else "10100" when (input = "00000000000100000000000000000000")
			else "10101" when (input = "00000000001000000000000000000000")
			else "10110" when (input = "00000000010000000000000000000000")
			else "10111" when (input = "00000000100000000000000000000000")
			else "11000" when (input = "00000001000000000000000000000000")
			else "11001" when (input = "00000010000000000000000000000000")
			else "11010" when (input = "00000100000000000000000000000000")
			else "11011" when (input = "00001000000000000000000000000000")
			else "11100" when (input = "00010000000000000000000000000000")
			else "11101" when (input = "00100000000000000000000000000000")
			else "11110" when (input = "01000000000000000000000000000000")
		   else "11111"; --when (input = "10000000000000000000000000000000");
		
			
end architecture behav;